`define BP_TWOBIT       (32'd0)
`define BP_GSHARE       (32'd1)
`define BP_GLOBAL       (32'd2)
`define BP_GSHARE_BASIC (32'd3)
`define BP_GLOBAL_BASIC (32'd4)
`define BP_LOCAL_BASIC  (32'd5)
`define BP_LOCAL_AHEAD  (32'd6)
`define BP_LOCAL_REPAIR (32'd7)